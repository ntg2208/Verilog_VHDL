module or_gate_code(a,b,y);

    input a,b;
    output y;
    
    assign y = a|b;

endmodule